LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY checker IS
  PORT (a_r: IN STD_LOGIC_VECTOR(22 DOWNTO 0);
        error: OUT STD_LOGIC);
END checker;

ARCHITECTURE Behavioral OF checker IS
BEGIN
END Behavioral;